module main

fn main() {
	println('learn quickjs tool')
}
